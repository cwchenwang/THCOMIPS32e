// Module RAMWrapper that adaptas SRAM modules as declared in thinpad_top.v 
// to a RAM module.
// With sel_i set to 4'b1111, this module can also be used to adapt SRAM to ROM.
// Author: LYL
// Created on: 2018/11/24

`timescale 1ns / 1ps
`include "defines.vh"

module RAMWrapper(
	input wire clk,
	
	// From MEM
    input wire ce_i,
    input wire we_i,
    input wire[`DataAddrBus] addr_i,
    input wire[3:0] sel_i,
    input wire[`DataBus] data_i,
    
    // To MEM
    output reg[`DataBus] data_o,
    
    // Adaptee
    inout wire[`InstBus] ram_data,  // RAM����
    output reg[19:0] ram_addr,      // RAM��ַ
    output reg[3:0] ram_be_n,       // RAM�ֽ�ʹ�ܣ�����Ч�������ʹ���ֽ�ʹ�ܣ��뱣��Ϊ0
    output reg ram_ce_n,            // RAMƬѡ������Ч
    output reg ram_oe_n,            // RAM��ʹ�ܣ�����Ч
    output reg ram_we_n             // RAMдʹ�ܣ�����Ч
);

    // Tri-state
    assign ram_data = (ce_i == `ChipEnable && we_i == `WriteEnable) ? data_i : {`DataWidth{1'bz}};
    
    // Read data_o from ram_data
    always @(*) begin
        if (ce_i == `ChipEnable && we_i == `WriteDisable) 
            data_o <= ram_data;
        else
            data_o <= 0;
    end
   
    always @ (*) begin
        ram_be_n <= 0;
        ram_addr <= addr_i[21:2];   // Only use low 20 bits, index by 32-bit word
        if (ce_i == `ChipDisable) begin
            ram_ce_n <= 1;
            ram_oe_n <= 1;
            ram_we_n <= 1;
        end else begin
            ram_ce_n <= 0;
            if (we_i == `WriteEnable) begin
                ram_oe_n <= 1;
                ram_we_n <= !clk;   // LOW at the first half cycle, HIGH for the rest
                ram_be_n <= ~sel_i;  // Happily, their meanings are almost the same
            end else begin  
                ram_oe_n <= 0;
                ram_we_n <= 1;
            end
        end
    end 
    
endmodule
